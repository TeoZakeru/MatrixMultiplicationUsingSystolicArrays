//module radix8_booth_multiplier #(parameter N = 8) (
//    input  signed [N-1:0] a,  // Multiplicand
//    input  signed [N-1:0] b,  // Multiplier
//    input clk, 
//    input rst,
//    output signed [2*N-1:0] Prod // Product
//);
//    localparam NUM_PARTIALS = (N + 2) / 3; // Compute ceil(N/3)	

//    reg signed [2*N:0] partial_products [NUM_PARTIALS-1:0]; // Array to store partial products
//    wire signed [2*N+1:0] accum; // Accumulator for final sum
//    wire [N+3:0] Q;
//    reg signed [3:0] booth_code [0:NUM_PARTIALS-1];
//    wire signed [N-1:0] neg_A;
//    wire signed [N:0] x2_A;
//    wire signed [N:0] x2_neg_A;
//    wire signed [N+1:0] x3_A;
//    wire signed [N+1:0] x3_neg_A;
//    wire signed [N+1:0] x4_A;
//    wire signed [N+1:0] x4_neg_A;
//    wire signed [N-1:0] A,B;
    
//    integer i;
//    always @(posedge clk or negedge rst) begin
//        if (!rst) begin
//            for (i = 0; i < NUM_PARTIALS; i = i + 1) begin
//                partial_products[i] <= 0;
//                booth_code[i] <= 0;
//            end
//        end else begin
//            for (i = 0; i < NUM_PARTIALS; i = i + 1) begin
//                booth_code[i] <= {Q[3*i+3], Q[3*i+2], Q[3*i+1], Q[3*i]};
//            end
//            for (i = 0; i < NUM_PARTIALS; i = i + 1) begin
//                case (booth_code[i])
//                    4'b0000, 4'b1111: partial_products[i] <= 0;
//                    4'b0001, 4'b0010: partial_products[i] <= {{(2*N+1-N){A[N-1]}}, A};       // +A
//                    4'b0011, 4'b0100: partial_products[i] <= {{(2*N+1-(N+1)){x2_A[N]}}, x2_A};  // +2A
//                    4'b0101, 4'b0110: partial_products[i] <= {{(2*N+1-(N+2)){x3_A[N+1]}}, x3_A}; // +3A
//                    4'b0111:          partial_products[i] <= {{(2*N+1-(N+2)){x4_A[N+1]}}, x4_A}; // +4A
//                    4'b1000:          partial_products[i] <= {{(2*N+1-(N+2)){x4_neg_A[N+1]}}, x4_neg_A}; // -4A
//                    4'b1001, 4'b1010: partial_products[i] <= {{(2*N+1-(N+2)){x3_neg_A[N+1]}}, x3_neg_A}; // -3A
//                    4'b1011, 4'b1100: partial_products[i] <= {{(2*N+1-(N+1)){x2_neg_A[N]}}, x2_neg_A};   // -2A
//                    4'b1101, 4'b1110: partial_products[i] <= {{(2*N+1-N){neg_A[N-1]}}, neg_A}; // -A
//                    default:          partial_products[i] <= 0;
//                endcase
//            end
//        end
//    end
    
//    assign accum = 
//        (partial_products[0] << (3*0)) +
//        (NUM_PARTIALS > 1 ? (partial_products[1] << (3*1)) : 0) +
//        (NUM_PARTIALS > 2 ? (partial_products[2] << (3*2)) : 0) +
//        (NUM_PARTIALS > 3 ? (partial_products[3] << (3*3)) : 0) +
//        (NUM_PARTIALS > 4 ? (partial_products[4] << (3*4)) : 0);
    
//    assign Q = {{3{B[N-1]}},B[N-1:0],1'b0};
//    assign A = (a[N-1] & b[N-1]) ? (~a + 1) : (b[N-1] ? b : a);
//    assign B = (a[N-1] & b[N-1]) ? (~b + 1) : (b[N-1] ? a : b);
//    // Compute 2's complement negation
//    assign neg_A = ~A + 1'b1;  
    
//    // Compute positive multiples with sign extension
//    assign x2_A = {A[N-1], A} << 1;  // 2A
//    assign x3_A = ({{2{A[N-1]}}, A} << 1) + {{2{A[N-1]}}, A}; // 3A = (2A + A)
//    assign x4_A = {{2{A[N-1]}}, A} << 2;  // 4A

//    // Compute negative multiples using 2's complement
//    assign x2_neg_A = (~{A[N-1], A} + 1'b1) << 1;  // -2A
//    assign x3_neg_A = {x2_neg_A[N-1],x2_neg_A} + {{2{neg_A[N-1]}},neg_A};// -3A
//    assign x4_neg_A = (~{{2{A[N-1]}}, A} + 1'b1) << 2;  // -4A
        
//    assign Prod = accum[2*N-1:0]; // Output the final product

//endmodule
module radix8_booth_multiplier #(parameter N = 8) (
    input  signed [N-1:0] a,  // Multiplicand
    input  signed [N-1:0] b,  // Multiplier
    input clk, 
    input rst,
    output reg [2*N-1:0] Prod // Product
);
    localparam NUM_PARTIALS = (N + 2) / 3; // Compute ceil(N/3)	
    reg signed [2*N:0] partial_products [NUM_PARTIALS-1:0]; // Array to store partial products
    wire signed [2*N+1:0] accum; // Accumulator for final sum
    wire [N+3:0] Q;
    wire signed [N-1:0] neg_A;
    wire signed [N:0] x2_A;
    wire signed [N:0] x2_neg_A;
    wire signed [N+1:0] x3_A;
    wire signed [N+1:0] x3_neg_A;
    wire signed [N+1:0] x4_A;
    wire signed [N+1:0] x4_neg_A;
    wire signed [N-1:0] A,B;
    reg signed [N-1:0] a_reg, b_reg;
    
    // Use generate for booth_code and partial_products logic
    integer i;
    wire [2*N-1:0] Product;
    
	always @(*) begin
        for (i = 0; i < NUM_PARTIALS; i = i + 1) begin : booth_encoding
                if (!rst) begin
                    partial_products[i] = 0;
                end else begin
                    case ({Q[3*i+3], Q[3*i+2], Q[3*i+1], Q[3*i]})
                        4'b0000, 4'b1111: partial_products[i] = 0;
                        4'b0001, 4'b0010: partial_products[i] = {{(2*N+1-N){A[N-1]}}, A};       // +A
                        4'b0011, 4'b0100: partial_products[i] = {{(2*N+1-(N+1)){x2_A[N]}}, x2_A};  // +2A
                        4'b0101, 4'b0110: partial_products[i] = {{(2*N+1-(N+2)){x3_A[N+1]}}, x3_A}; // +3A
                        4'b0111:          partial_products[i] = {{(2*N+1-(N+2)){x4_A[N+1]}}, x4_A}; // +4A
                        4'b1000:          partial_products[i] = {{(2*N+1-(N+2)){x4_neg_A[N+1]}}, x4_neg_A}; // -4A
                        4'b1001, 4'b1010: partial_products[i] = {{(2*N+1-(N+2)){x3_neg_A[N+1]}}, x3_neg_A}; // -3A
                        4'b1011, 4'b1100: partial_products[i] = {{(2*N+1-(N+1)){x2_neg_A[N]}}, x2_neg_A};   // -2A
                        4'b1101, 4'b1110: partial_products[i] = {{(2*N+1-N){neg_A[N-1]}}, neg_A}; // -A
                        default:          partial_products[i] = 0;
                    endcase
                end
            end
        end
    
    // Accumulate partial products using generate
//    generate
//        if (NUM_PARTIALS == 1) begin : single_partial
//            assign accum = partial_products[0] << (3*0);
//        end else if (NUM_PARTIALS == 2) begin : two_partials
//            assign accum = (partial_products[0] << (3*0)) +
//                           (partial_products[1] << (3*1));
//        end else if (NUM_PARTIALS == 3) begin : three_partials
//            assign accum = (partial_products[0] << (3*0)) +
//                           (partial_products[1] << (3*1)) +
//                           (partial_products[2] << (3*2));
//        end else if (NUM_PARTIALS == 4) begin : four_partials
//            assign accum = (partial_products[0] << (3*0)) +
//                           (partial_products[1] << (3*1)) +
//                           (partial_products[2] << (3*2)) +
//                           (partial_products[3] << (3*3));
//        end else begin : five_plus_partials
//            assign accum = (partial_products[0] << (3*0)) +
//                           (partial_products[1] << (3*1)) +
//                           (partial_products[2] << (3*2)) +
//                           (partial_products[3] << (3*3)) +
//                           (partial_products[4] << (3*4));
//        end
//    endgenerate

	always @(posedge clk or negedge rst) begin
		if(!rst) begin
			a_reg <= 0;
			b_reg <= 0;
			Prod <= 0;
		end
		else begin
			a_reg <= a;
			b_reg <= b;
			Prod <= Product;
		end
	end

	WallaceTreeMult mul(
		.clk(clk),
		.rst(rst),
		.P1_in(partial_products[0][31:0]),
		.P2_in(partial_products[1][28:0]),
		.P3_in(partial_products[2][25:0]),
		.P4_in(partial_products[3][22:0]),
		.P5_in(partial_products[4][19:0]),
		.P6_in(partial_products[5][16:0]),
		.Out(Product)
    );
    
    assign Q = {{3{B[N-1]}},B[N-1:0],1'b0};
    assign A = (a_reg[N-1] & b_reg[N-1]) ? (~a_reg + 1) : (b_reg[N-1] ? b_reg : a_reg);
    assign B = (a_reg[N-1] & b_reg[N-1]) ? (~b_reg + 1) : (b_reg[N-1] ? a_reg : b_reg);
    // Compute 2's complement negation
    assign neg_A = ~A + 1'b1;  
    
    // Compute positive multiples with sign extension
    assign x2_A = {A[N-1], A} << 1;  // 2A
    assign x3_A = ({{2{A[N-1]}}, A} << 1) + {{2{A[N-1]}}, A}; // 3A = (2A + A)
    assign x4_A = {{2{A[N-1]}}, A} << 2;  // 4A
    // Compute negative multiples using 2's complement
    assign x2_neg_A = (~{A[N-1], A} + 1'b1) << 1;  // -2A
    assign x3_neg_A = {x2_neg_A[N-1],x2_neg_A} + {{2{neg_A[N-1]}},neg_A};// -3A
    assign x4_neg_A = (~{{2{A[N-1]}}, A} + 1'b1) << 2;  // -4A
        
//    assign Prod = accum[2*N-1:0]; // Output the final product
endmodule
