`timescale 1ns / 1ps

module SA_tb;

    parameter SIZE = 8;
    parameter DATA_WIDTH = 16;

    // Inputs
    reg clk;
    reg rst;
    reg [SIZE*DATA_WIDTH-1:0] A;
    reg [SIZE*DATA_WIDTH-1:0] B;
    wire [SIZE*SIZE*2*DATA_WIDTH-1:0] C;
    // Outputs
    wire done;
    // Instantiate the SA module
    SystolicArray #(.SIZE(SIZE), .DATA_WIDTH(DATA_WIDTH)) uut (
        .A(A),
        .B(B),
        .clk(clk),
        .rst(rst),
        .done(done),
        .C(C)
    );

    // Clock generation (50% duty cycle, period = 10ns)
    always #5 clk = ~clk;
    initial begin
    $dumpfile("wave.vcd");
    $dumpvars(0, SA_tb);
    end

    initial begin
        #150;
        clk = 0;
        rst = 0;
        #10 rst = 1;
        $monitor("%t %h", $time, C);

        A = {16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd37};
        B = {16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd2};
        #10;
        A = {16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd45, 16'd60};
        B = {16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd30, 16'd47};
        #10;
        A = {16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd53, 16'd45, 16'd1};
        B = {16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd27, 16'd25, 16'd2};
        #10;
        A = {16'd0, 16'd0, 16'd0, 16'd0, 16'd49, 16'd63, 16'd40, 16'd5};
        B = {16'd0, 16'd0, 16'd0, 16'd0, 16'd48, 16'd61, 16'd56, 16'd5};
        #10;
        A = {16'd0, 16'd0, 16'd0, 16'd14, 16'd24, 16'd35, 16'd48, 16'd52};
        B = {16'd0, 16'd0, 16'd0, 16'd2, 16'd57, 16'd1, 16'd46, 16'd16};
        #10;
        A = {16'd0, 16'd0, 16'd61, 16'd50, 16'd7, 16'd31, 16'd23, 16'd23};
        B = {16'd0, 16'd0, 16'd57, 16'd11, 16'd45, 16'd22, 16'd4, 16'd48};
        #10;
        A = {16'd0, 16'd0, 16'd3, 16'd53, 16'd28, 16'd19, 16'd12, 16'd44};
        B = {16'd0, 16'd42, 16'd22, 16'd42, 16'd2, 16'd19, 16'd23, 16'd46};
        #10;
        A = {16'd56, 16'd46, 16'd54, 16'd56, 16'd38, 16'd35, 16'd29, 16'd50};
        B = {16'd6, 16'd14, 16'd32, 16'd5, 16'd39, 16'd48, 16'd4, 16'd53};
        #10;
        A = {16'd56, 16'd1, 16'd22, 16'd53, 16'd59, 16'd59, 16'd50, 16'd0};
        B = {16'd56, 16'd52, 16'd17, 16'd28, 16'd54, 16'd38, 16'd8, 16'd0};
        #10;
        A = {16'd7, 16'd32, 16'd28, 16'd58, 16'd7, 16'd62, 16'd0, 16'd0};
        B = {16'd56, 16'd2, 16'd0, 16'd7, 16'd15, 16'd47, 16'd0, 16'd0};
        #10;
        A = {16'd42, 16'd9, 16'd13, 16'd19, 16'd19, 16'd0, 16'd0, 16'd0};
        B = {16'd12, 16'd58, 16'd2, 16'd60, 16'd5, 16'd0, 16'd0, 16'd0};
        #10;
        A = {16'd51, 16'd51, 16'd27, 16'd21, 16'd0, 16'd0, 16'd0, 16'd0};
        B = {16'd60, 16'd48, 16'd11, 16'd31, 16'd0, 16'd0, 16'd0, 16'd0};
        #10;
        A = {16'd35, 16'd17, 16'd33, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0};
        B = {16'd51, 16'd1, 16'd16, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0};
        #10;
        A = {16'd3, 16'd62, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0};
        B = {16'd28, 16'd18, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0};
        #10;
        A = {16'd13, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0};
        B = {16'd40, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0};
        #10;
        A = 128'd0;
        B = 128'd0;
        #10;
        A = 128'd0;
        B = 128'd0;
        #10;
        A = 128'd0;
        B = 128'd0;
        #10;
        A = 128'd0;
        B = 128'd0;
        #10;
        A = 128'd0;
        B = 128'd0;
        #10;
        A = 128'd0;
        B = 128'd0;
        #10;
        A = 128'd0;
        B = 128'd0;
        #10;
        A = 128'd0;
        B = 128'd0;

    end
    
    endmodule

