`timescale 1ns / 1ps

module SA_tb;

    parameter SIZE = 8;
    parameter DATA_WIDTH = 32;

    // Inputs
    reg clk;
    reg rst;
    reg [SIZE*DATA_WIDTH-1:0] A;
    reg [SIZE*DATA_WIDTH-1:0] B;
    wire [SIZE*SIZE*2*DATA_WIDTH-1:0] C;
    // Outputs
    wire done;
    // Instantiate the SA module
    SystolicArray #(.SIZE(SIZE), .DATA_WIDTH(DATA_WIDTH)) uut (
        .A(A),
        .B(B),
        .clk(clk),
        .rst(rst),
        .done(done),
        .C(C)
    );

    // Clock generation (50% duty cycle, period = 10ns)
    always #5 clk = ~clk;
    initial begin
    $dumpfile("wave.vcd");
    $dumpvars(0, SA_tb);
    end

    initial begin
        #150;
        clk = 0;
        rst = 0;
        #10 rst = 1;
        $monitor("%t %h", $time, C);

        A = {32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd37};
        B = {32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd2};
        #10;
        A = {32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd45, 32'd60};
        B = {32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd30, 32'd47};
        #10;
        A = {32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd53, 32'd45, 32'd1};
        B = {32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd27, 32'd25, 32'd2};
        #10;
        A = {32'd0, 32'd0, 32'd0, 32'd0, 32'd49, 32'd63, 32'd40, 32'd5};
        B = {32'd0, 32'd0, 32'd0, 32'd0, 32'd48, 32'd61, 32'd56, 32'd5};
        #10;
        A = {32'd0, 32'd0, 32'd0, 32'd14, 32'd24, 32'd35, 32'd48, 32'd52};
        B = {32'd0, 32'd0, 32'd0, 32'd2, 32'd57, 32'd1, 32'd46, 32'd16};
        #10;
        A = {32'd0, 32'd0, 32'd61, 32'd50, 32'd7, 32'd31, 32'd23, 32'd23};
        B = {32'd0, 32'd0, 32'd57, 32'd11, 32'd45, 32'd22, 32'd4, 32'd48};
        #10;
        A = {32'd0, 32'd0, 32'd3, 32'd53, 32'd28, 32'd19, 32'd12, 32'd44};
        B = {32'd0, 32'd42, 32'd22, 32'd42, 32'd2, 32'd19, 32'd23, 32'd46};
        #10;
        A = {32'd56, 32'd46, 32'd54, 32'd56, 32'd38, 32'd35, 32'd29, 32'd50};
        B = {32'd6, 32'd14, 32'd32, 32'd5, 32'd39, 32'd48, 32'd4, 32'd53};
        #10;
        A = {32'd56, 32'd1, 32'd22, 32'd53, 32'd59, 32'd59, 32'd50, 32'd0};
        B = {32'd56, 32'd52, 32'd17, 32'd28, 32'd54, 32'd38, 32'd8, 32'd0};
        #10;
        A = {32'd7, 32'd32, 32'd28, 32'd58, 32'd7, 32'd62, 32'd0, 32'd0};
        B = {32'd56, 32'd2, 32'd0, 32'd7, 32'd15, 32'd47, 32'd0, 32'd0};
        #10;
        A = {32'd42, 32'd9, 32'd13, 32'd19, 32'd19, 32'd0, 32'd0, 32'd0};
        B = {32'd12, 32'd58, 32'd2, 32'd60, 32'd5, 32'd0, 32'd0, 32'd0};
        #10;
        A = {32'd51, 32'd51, 32'd27, 32'd21, 32'd0, 32'd0, 32'd0, 32'd0};
        B = {32'd60, 32'd48, 32'd11, 32'd31, 32'd0, 32'd0, 32'd0, 32'd0};
        #10;
        A = {32'd35, 32'd17, 32'd33, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0};
        B = {32'd51, 32'd1, 32'd16, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0};
        #10;
        A = {32'd3, 32'd62, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0};
        B = {32'd28, 32'd18, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0};
        #10;
        A = {32'd13, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0};
        B = {32'd40, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0};
        #10;
        A = 256'd0;
        B = 256'd0;
        #10;
        A = 256'd0;
        B = 256'd0;
        #10;
        A = 256'd0;
        B = 256'd0;
        #10;
        A = 256'd0;
        B = 256'd0;
        #10;
        A = 256'd0;
        B = 256'd0;
        #10;
        A = 256'd0;
        B = 256'd0;
        #10;
        A = 256'd0;
        B = 256'd0;
        #10;
        A = 256'd0;
        B = 256'd0;

    end
    
    endmodule

