//`timescale 1ns / 1ps

//module SA_tb;

//    parameter SIZE = 2;
//    parameter DATA_WIDTH = 8;

//    // Inputs
//    reg clk;
//    reg rst;
//    reg [SIZE*DATA_WIDTH-1:0] A;
//    reg [SIZE*DATA_WIDTH-1:0] B;
//    wire [SIZE*SIZE*2*DATA_WIDTH-1:0] C;
//    reg start;
//    // Outputs
//    wire done;
//    // Instantiate the SA module
//    SystolicArray #(.SIZE(SIZE), .DATA_WIDTH(DATA_WIDTH)) uut (
//        .A(A),
//        .B(B),
//        .clk(clk),
//        .rst(rst),
//        .done(done),
//        .C(C),
//        .start(start)
//    );

//    // Clock generation (50% duty cycle, period = 10ns)
//    always #5 clk = ~clk;

//    // Task to print the output matrix

//    // Test procedure
//    initial begin
//    	#150;
//		clk = 0;
//		start = 0;
//        // Initialize clock and reset
//        rst = 0;
//		#100;
//        #10 rst = 1; // Release reset after 10ns
//        // Initialize input matrices A and B (row-major order)
//        start = 1'b1;
//        A = {8'd0, 8'd1};
//        B = {8'd0, 8'd4};
//        #10;
//        A = {8'd3, 8'd2};
//        B = {8'd3, 8'd2};
//        #10;
//        A = {8'd4, 8'd0};
//        B = {8'd1, 8'd0};
////        #10;
////        A = {8'd0, 8'd0};
////        B = {8'd0, 8'd0};
////        #10;
////        A = {8'd0, 8'd0};
////        B = {8'd0, 8'd0};
//        #10;
//        A = {8'd0, 8'd5};
//        B = {8'd0, 8'd1};;
//        #10;
//        A = {8'd7, 8'd6};
//        B = {8'd3, 8'd2};
//        #10;
//        A = {8'd8, 8'd0};
//        B = {8'd4, 8'd0};
//        #10;
//        A = {8'd0, 8'd0};
//        B = {8'd0, 8'd0};
//        #10;
//        A = {8'd0, 8'd0};
//        B = {8'd0, 8'd0};
//        #10;
//        A = {8'd0, 8'd0};
//        B = {8'd0, 8'd0};
////		A = {9'd0,9'd0,9'd4};
////		B = {9'd0,9'd0,9'd6};
////		#10;
////		A = {9'd0,9'd16,9'd5};
////		B = {9'd0,9'd12,9'd19};
////		#10;
////		A = {9'd2,9'd5,9'd7};
////		B = {9'd2,9'd7,9'd18};
////		#10;
////		A = {9'd8,9'd15,9'd0};
////		B = {9'd16,9'd2,9'd0};
////		#10;
////		A = {9'd4,9'd0,9'd0};
////		B = {9'd18,9'd0,9'd0};
////		#10;
////		A = {9'd0,9'd0,9'd0};
////		B = {9'd0,9'd0,9'd0};
////		#10;
////		A = {9'd0,9'd0,9'd0};
////		B = {9'd0,9'd0,9'd0};
////		#10;A = {9'd0,9'd0,9'd0};
////		B = {9'd0,9'd0,9'd0};
////		#10;
////		A = {9'd0,9'd0,9'd0};
////		B = {9'd0,9'd0,9'd0};
////		#10;A = {9'd0,9'd0,9'd0};
////		B = {9'd0,9'd0,9'd0};
////		#10;
////		A = {9'd0,9'd0,9'd0};
////		B = {9'd0,9'd0,9'd0};
////		#10;
		
//        // Wait for computation to complete
//        wait(done);

//        // Print output matrix
//        #1000;
//    end
//endmodule


`timescale 1ns / 1ps

module SA_tb;

    parameter SIZE = 8;
    parameter DATA_WIDTH = 8;

    // Inputs
    reg clk;
    reg rst;
    reg [SIZE*DATA_WIDTH-1:0] A;
    reg [SIZE*DATA_WIDTH-1:0] B;
    wire [SIZE*SIZE*2*DATA_WIDTH-1:0] C;
    // Outputs
    wire done;
    reg start;
    // Instantiate the SA module
    SystolicArray #(.SIZE(SIZE), .DATA_WIDTH(DATA_WIDTH)) uut (
        .A(A),
        .B(B),
        .clk(clk),
        .rst(rst),
        .done(done),
        .C(C),
        .start(start)
    );

    // Clock generation (50% duty cycle, period = 10ns)
    always #5 clk = ~clk;

    // Task to print the output matrix

    // Test procedure
//    initial begin
//    $dumpfile("wave.vcd");
//    $dumpvars(0, SA_tb);
//    end 
//    initial begin
//    	#150;
//		clk = 0;
//        // Initialize clock and reset
//        rst = 0;
//        #10 rst = 1; // Release reset after 10ns
//        // Initialize input matrices A and B (row-major order)
        

////8x8 matrix

//    A = {8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd1};
//    B = {8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd1};
//    #10;
//    A = {8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd2, 8'd1};
//    B = {8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd2, 8'd1};
//    #10;
//    A = {8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd3, 8'd2, 8'd1};
//    B = {8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd3, 8'd2, 8'd1};
//    #10;
//    A = {8'd0, 8'd0, 8'd0, 8'd0, 8'd4, 8'd3, 8'd2, 8'd1};
//    B = {8'd0, 8'd0, 8'd0, 8'd0, 8'd4, 8'd3, 8'd2, 8'd1};
//    #10;
//    A = {8'd0, 8'd0, 8'd0, 8'd5, 8'd4, 8'd3, 8'd2, 8'd1};
//    B = {8'd0, 8'd0, 8'd0, 8'd5, 8'd4, 8'd3, 8'd2, 8'd1};
//    #10;
//    A = {8'd0, 8'd0, 8'd6, 8'd5, 8'd4, 8'd3, 8'd2, 8'd1};
//    B = {8'd0, 8'd0, 8'd6, 8'd5, 8'd4, 8'd3, 8'd2, 8'd1};
//    #10;
//    A = {8'd0, 8'd7, 8'd6, 8'd5, 8'd4, 8'd3, 8'd2, 8'd1};
//    B = {8'd0, 8'd7, 8'd6, 8'd5, 8'd4, 8'd3, 8'd2, 8'd1};
//    #10;
//    A = {8'd8, 8'd7, 8'd6, 8'd5, 8'd4, 8'd3, 8'd2, 8'd1};
//    B = {8'd8, 8'd7, 8'd6, 8'd5, 8'd4, 8'd3, 8'd2, 8'd1};        
//	#10;
//    A = {8'd8, 8'd7, 8'd6, 8'd5, 8'd4, 8'd3, 8'd2, 8'd0};
//    B = {8'd8, 8'd7, 8'd6, 8'd5, 8'd4, 8'd3, 8'd2, 8'd0}; 
//	#10;
//    A = {8'd8, 8'd7, 8'd6, 8'd5, 8'd4, 8'd3, 8'd0, 8'd0};
//    B = {8'd8, 8'd7, 8'd6, 8'd5, 8'd4, 8'd3, 8'd0, 8'd0};
//	#10;
//    A = {8'd8, 8'd7, 8'd6, 8'd5, 8'd4, 8'd0, 8'd0, 8'd0};
//    B = {8'd8, 8'd7, 8'd6, 8'd5, 8'd4, 8'd0, 8'd0, 8'd0};
//    #10;
//    A = {8'd8, 8'd7, 8'd6, 8'd5, 8'd0, 8'd0, 8'd0, 8'd0};
//    B = {8'd8, 8'd7, 8'd6, 8'd5, 8'd0, 8'd0, 8'd0, 8'd0};
//    #10;
//    A = {8'd8, 8'd7, 8'd6, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0};
//    B = {8'd8, 8'd7, 8'd6, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0};
//    #10;
//    A = {8'd8, 8'd7, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0};
//    B = {8'd8, 8'd7, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0};
//    #10;
//    A = {8'd8, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0};
//    B = {8'd8, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0};
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
//	A = 64'd0;
//	B = 64'd0;
//	#10;
	

//        // Wait for computation to complete
//    wait(done);

//        // Print output matrix
//        // $displ
////        #1000;
//        #60;        
//        // End simulation
//        $stop;
//    end
//endmodule
wire [2*DATA_WIDTH-1:0] C_unpacked [0:SIZE-1][0:SIZE-1];
		genvar i, j;
generate
    for (i = 0; i < SIZE; i = i + 1) begin : row_loop
        for (j = 0; j < SIZE; j = j + 1) begin : col_loop
            assign C_unpacked[i][j] = C[(i*SIZE + j + 1)*2*DATA_WIDTH - 1 -: 2*DATA_WIDTH];
        end
    end
endgenerate

    initial begin
    $dumpfile("wave.vcd");
    $dumpvars(0, SA_tb);
    end

    initial begin
    	$monitor("%t %h",$time, C);
        #150;
        clk = 0;
        rst = 0;
        #10 rst = 1;
//        #5;
		start = 1;
       	A  = {8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd37};
        B = {8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd2};
        #10;
        A = {8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd45, 8'd60};
        B = {8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd30, 8'd47};
        #10;
        A = {8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd53, 8'd45, 8'd1};
        B = {8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd27, 8'd25, 8'd2};
        #10;
        A = {8'd0, 8'd0, 8'd0, 8'd0, 8'd49, 8'd63, 8'd40, 8'd5};
        B = {8'd0, 8'd0, 8'd0, 8'd0, 8'd48, 8'd61, 8'd56, 8'd5};
        #10;
        A = {8'd0, 8'd0, 8'd0, 8'd14, 8'd24, 8'd35, 8'd48, 8'd52};
        B = {8'd0, 8'd0, 8'd0, 8'd2, 8'd57, 8'd1, 8'd46, 8'd16};
        #10;
        A = {8'd0, 8'd0, 8'd61, 8'd50, 8'd7, 8'd31, 8'd23, 8'd23};
        B = {8'd0, 8'd0, 8'd57, 8'd11, 8'd45, 8'd22, 8'd4, 8'd48};
        #10;
        A = {8'd0, 8'd0, 8'd3, 8'd53, 8'd28, 8'd19, 8'd12, 8'd44};
        B = {8'd0, 8'd42, 8'd22, 8'd42, 8'd2, 8'd19, 8'd23, 8'd46};
        #10;
        A = {8'd56, 8'd46, 8'd54, 8'd56, 8'd38, 8'd35, 8'd29, 8'd50};
        B = {8'd6, 8'd14, 8'd32, 8'd5, 8'd39, 8'd48, 8'd4, 8'd53};
        #10;
        A = {8'd56, 8'd1, 8'd22, 8'd53, 8'd59, 8'd59, 8'd50, 8'd0};
        B = {8'd56, 8'd52, 8'd17, 8'd28, 8'd54, 8'd38, 8'd8, 8'd0};
        #10;
        A = {8'd7, 8'd32, 8'd28, 8'd58, 8'd7, 8'd62, 8'd0, 8'd0};
        B = {8'd56, 8'd2, 8'd0, 8'd7, 8'd15, 8'd47, 8'd0, 8'd0};
        #10;
        A = {8'd42, 8'd9, 8'd13, 8'd19, 8'd19, 8'd0, 8'd0, 8'd0};
        B = {8'd12, 8'd58, 8'd2, 8'd60, 8'd5, 8'd0, 8'd0, 8'd0};
        #10;
        A = {8'd51, 8'd51, 8'd27, 8'd21, 8'd0, 8'd0, 8'd0, 8'd0};
        B = {8'd60, 8'd48, 8'd11, 8'd31, 8'd0, 8'd0, 8'd0, 8'd0};
        #10;
        A = {8'd35, 8'd17, 8'd33, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0};
        B = {8'd51, 8'd1, 8'd16, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0};
        #10;
        A = {8'd3, 8'd62, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0};
        B = {8'd28, 8'd18, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0};
        #10;
        A = {8'd13, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0};
        B = {8'd40, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0};
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;
        A  = {8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd37};
        B = {8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd2};
        #10;
        A = {8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd45, 8'd60};
        B = {8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd30, 8'd47};
        #10;
        A = {8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd53, 8'd45, 8'd1};
        B = {8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd27, 8'd25, 8'd2};
        #10;
        A = {8'd0, 8'd0, 8'd0, 8'd0, 8'd49, 8'd63, 8'd40, 8'd5};
        B = {8'd0, 8'd0, 8'd0, 8'd0, 8'd48, 8'd61, 8'd56, 8'd5};
        #10;
        A = {8'd0, 8'd0, 8'd0, 8'd14, 8'd24, 8'd35, 8'd48, 8'd52};
        B = {8'd0, 8'd0, 8'd0, 8'd2, 8'd57, 8'd1, 8'd46, 8'd16};
        #10;
        A = {8'd0, 8'd0, 8'd61, 8'd50, 8'd7, 8'd31, 8'd23, 8'd23};
        B = {8'd0, 8'd0, 8'd57, 8'd11, 8'd45, 8'd22, 8'd4, 8'd48};
        #10;
        A = {8'd0, 8'd0, 8'd3, 8'd53, 8'd28, 8'd19, 8'd12, 8'd44};
        B = {8'd0, 8'd42, 8'd22, 8'd42, 8'd2, 8'd19, 8'd23, 8'd46};
        #10;
        A = {8'd56, 8'd46, 8'd54, 8'd56, 8'd38, 8'd35, 8'd29, 8'd50};
        B = {8'd6, 8'd14, 8'd32, 8'd5, 8'd39, 8'd48, 8'd4, 8'd53};
        #10;
        A = {8'd56, 8'd1, 8'd22, 8'd53, 8'd59, 8'd59, 8'd50, 8'd0};
        B = {8'd56, 8'd52, 8'd17, 8'd28, 8'd54, 8'd38, 8'd8, 8'd0};
        #10;
        A = {8'd7, 8'd32, 8'd28, 8'd58, 8'd7, 8'd62, 8'd0, 8'd0};
        B = {8'd56, 8'd2, 8'd0, 8'd7, 8'd15, 8'd47, 8'd0, 8'd0};
        #10;
        A = {8'd42, 8'd9, 8'd13, 8'd19, 8'd19, 8'd0, 8'd0, 8'd0};
        B = {8'd12, 8'd58, 8'd2, 8'd60, 8'd5, 8'd0, 8'd0, 8'd0};
        #10;
        A = {8'd51, 8'd51, 8'd27, 8'd21, 8'd0, 8'd0, 8'd0, 8'd0};
        B = {8'd60, 8'd48, 8'd11, 8'd31, 8'd0, 8'd0, 8'd0, 8'd0};
        #10;
        A = {8'd35, 8'd17, 8'd33, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0};
        B = {8'd51, 8'd1, 8'd16, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0};
        #10;
        A = {8'd3, 8'd62, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0};
        B = {8'd28, 8'd18, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0};
        #10;
        A = {8'd13, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0};
        B = {8'd40, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0};
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;
        A = 64'd0;
        B = 64'd0;
        #10;

        wait(done);
        #60;
        #10000;
        
    end
    
    endmodule
